class AXI_M_w_monitor extends uvm_monitor;

  `uvm_component_utils(AXI_M_w_monitor)
  
  // declaring virual interface
  virtual interface AXI4_if vif;

  // Collected Data handle
  AXI_M_w_txn pkt;

  // Count packets collected
  int num_pkt_col;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("Monitor", "Inside AXI_M_w_monitor build_phase", UVM_LOW)
  endfunction

  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    if (!uvm_config_db#(virtual AXI4_if)::get(this, "", "vif", vif)) begin
      `uvm_fatal(get_type_name(), "NO-VIF")
    end
  endfunction

  task run_phase(uvm_phase phase);
    `uvm_info("Monitor", "Inside AXI_M_w_monitor run_phase", UVM_LOW)
    monitor_write();
  endtask

  task monitor_write();
    forever begin
      // Wait for reset deassertion
      @(posedge vif.ACLK);
      wait(vif.ARESETn == 1);

      // Wait for AWVALID and AWREADY handshake
      if (vif.AWVALID && vif.AWREADY) begin
        pkt = AXI_M_w_txn::type_id::create("pkt");
        pkt.AWADDR  = vif.AWADDR;
        pkt.AWVALID = vif.AWVALID;
        pkt.AWREADY = vif.AWREADY;

        // Wait for WVALID and WREADY handshake
        if (vif.WVALID && vif.WREADY) begin
          pkt.WDATA  = vif.WDATA;
          pkt.WVALID = vif.WVALID;
          pkt.WREADY = vif.WREADY;

          num_pkt_col++;
          `uvm_info("Monitor", $sformatf("Collected Write txn %0d: AWADDR=0x%0h WDATA=0x%0h", num_pkt_col, pkt.AWADDR, pkt.WDATA), UVM_LOW);
        end
      end
    end
  endtask
endclass
